/**
  @brief A module of mysterious purpose

  @input clk    clock
  @input nReset active-low reset
  @input a      an input
  @input b      an input
  @input c      an input

  @output out   output
*/
module Exercise3 (
    input clk,
    input nReset,
    input [3:0] a,
    input [15:0] b,
    input [15:0] c,
    output [15:0] out
);

endmodule
